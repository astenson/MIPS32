/*******************************************************************************
Project: 32-bit Out of Order MIPS Processor
Author: Adam Stenson
Module: MIPS, overall pipeline connecting individual component blocks
Last Updated: December 21, 2018
*******************************************************************************/

module MIPS();

endmodule
